module FFT_Processor();

endmodule