module clkdiv50to4_TB;

	reg clk50;
	wire clk4;
	
	clkdiv50to4 UUT(clk50, clk4);
	
	initial begin
		clk50 = 1;
		#10;
		clk50 = 0;
		#10;
		clk50 = 1;
		#10;
		clk50 = 0;
		#10;
		clk50 = 1;
		#10;
		clk50 = 0;
		#10;
		clk50 = 1;
		#10;
		clk50 = 0;
		#10;
		clk50 = 1;
		#10;
		clk50 = 0;
		#10;
		clk50 = 1;
		#10;
		clk50 = 0;
		#10;
		clk50 = 1;
		#10;
		clk50 = 0;
		#10;
		clk50 = 1;
		#10;
		clk50 = 0;
		#10;
		clk50 = 1;
		#10;
		clk50 = 0;
		#10;
		clk50 = 1;
		#10;
		clk50 = 0;
		#10;
		clk50 = 1;
		#10;
		clk50 = 0;
		#10;
		clk50 = 1;
		#10;
		clk50 = 0;
		#10;
		clk50 = 1;
		#10;
		clk50 = 0;
		#10;
		clk50 = 1;
		#10;
		clk50 = 0;
		#10;
		clk50 = 1;
		#10;
		clk50 = 0;
		#10;
		clk50 = 1;
		#10;
		clk50 = 0;
		#10;
		clk50 = 1;
		#10;
		clk50 = 0;
		#10;
		clk50 = 1;
		#10;
		clk50 = 0;
		#10;
	end

endmodule